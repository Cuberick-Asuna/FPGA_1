module f2_ROM ( input wire [3:0] x,
input wire [3:0] y,
input wire [1:0] image_no,
output wire [2:0] color
);

reg [2:0] current_pxl_color;
wire [7:0] pxl_coor;

assign pxl_coor = {x,y};


always @(*)
begin
	case (image_no)
		0  :
			begin
				case (pxl_coor)
					0	: current_pxl_color = 3'b111;
					1	: current_pxl_color = 3'b111;
					2	: current_pxl_color = 3'b111;
					3	: current_pxl_color = 3'b111;
					4	: current_pxl_color = 3'b111;
					5	: current_pxl_color = 3'b111;
					6	: current_pxl_color = 3'b111;
					7	: current_pxl_color = 3'b111;
					8	: current_pxl_color = 3'b111;
					9	: current_pxl_color = 3'b111;
					10	: current_pxl_color = 3'b111;
					11	: current_pxl_color = 3'b111;
					12	: current_pxl_color = 3'b111;
					13	: current_pxl_color = 3'b111;
					14	: current_pxl_color = 3'b111;
					15	: current_pxl_color = 3'b111;
					16	: current_pxl_color = 3'b111;
					17	: current_pxl_color = 3'b111;
					18	: current_pxl_color = 3'b111;
					19	: current_pxl_color = 3'b111;
					20	: current_pxl_color = 3'b111;
					21	: current_pxl_color = 3'b111;
					22	: current_pxl_color = 3'b000;
					23	: current_pxl_color = 3'b000;
					24	: current_pxl_color = 3'b000;
					25	: current_pxl_color = 3'b000;
					26	: current_pxl_color = 3'b111;
					27	: current_pxl_color = 3'b111;
					28	: current_pxl_color = 3'b111;
					29	: current_pxl_color = 3'b111;
					30	: current_pxl_color = 3'b111;
					31	: current_pxl_color = 3'b111;
					32	: current_pxl_color = 3'b111;
					33	: current_pxl_color = 3'b111;
					34	: current_pxl_color = 3'b111;
					35	: current_pxl_color = 3'b111;
					36	: current_pxl_color = 3'b111;
					37	: current_pxl_color = 3'b000;
					38	: current_pxl_color = 3'b000;
					39	: current_pxl_color = 3'b000;
					40	: current_pxl_color = 3'b000;
					41	: current_pxl_color = 3'b000;
					42	: current_pxl_color = 3'b000;
					43	: current_pxl_color = 3'b111;
					44	: current_pxl_color = 3'b111;
					45	: current_pxl_color = 3'b111;
					46	: current_pxl_color = 3'b111;
					47	: current_pxl_color = 3'b111;
					48	: current_pxl_color = 3'b111;
					49	: current_pxl_color = 3'b111;
					50	: current_pxl_color = 3'b111;
					51	: current_pxl_color = 3'b111;
					52	: current_pxl_color = 3'b000;
					53	: current_pxl_color = 3'b000;
					54	: current_pxl_color = 3'b111;
					55	: current_pxl_color = 3'b111;
					56	: current_pxl_color = 3'b111;
					57	: current_pxl_color = 3'b111;
					58	: current_pxl_color = 3'b000;
					59	: current_pxl_color = 3'b000;
					60	: current_pxl_color = 3'b111;
					61	: current_pxl_color = 3'b111;
					62	: current_pxl_color = 3'b111;
					63	: current_pxl_color = 3'b111;
					64	: current_pxl_color = 3'b111;
					65	: current_pxl_color = 3'b111;
					66	: current_pxl_color = 3'b111;
					67	: current_pxl_color = 3'b111;
					68	: current_pxl_color = 3'b000;
					69	: current_pxl_color = 3'b111;
					70	: current_pxl_color = 3'b111;
					71	: current_pxl_color = 3'b111;
					72	: current_pxl_color = 3'b111;
					73	: current_pxl_color = 3'b111;
					74	: current_pxl_color = 3'b111;
					75	: current_pxl_color = 3'b000;
					76	: current_pxl_color = 3'b111;
					77	: current_pxl_color = 3'b111;
					78	: current_pxl_color = 3'b111;
					79	: current_pxl_color = 3'b111;
					80	: current_pxl_color = 3'b111;
					81	: current_pxl_color = 3'b111;
					82	: current_pxl_color = 3'b111;
					83	: current_pxl_color = 3'b111;
					84	: current_pxl_color = 3'b000;
					85	: current_pxl_color = 3'b111;
					86	: current_pxl_color = 3'b000;
					87	: current_pxl_color = 3'b111;
					88	: current_pxl_color = 3'b111;
					89	: current_pxl_color = 3'b000;
					90	: current_pxl_color = 3'b111;
					91	: current_pxl_color = 3'b000;
					92	: current_pxl_color = 3'b111;
					93	: current_pxl_color = 3'b111;
					94	: current_pxl_color = 3'b111;
					95	: current_pxl_color = 3'b111;
					96	: current_pxl_color = 3'b111;
					97	: current_pxl_color = 3'b111;
					98	: current_pxl_color = 3'b111;
					99	: current_pxl_color = 3'b000;
					100	: current_pxl_color = 3'b000;
					101	: current_pxl_color = 3'b111;
					102	: current_pxl_color = 3'b000;
					103	: current_pxl_color = 3'b111;
					104	: current_pxl_color = 3'b111;
					105	: current_pxl_color = 3'b000;
					106	: current_pxl_color = 3'b111;
					107	: current_pxl_color = 3'b000;
					108	: current_pxl_color = 3'b000;
					109	: current_pxl_color = 3'b111;
					110	: current_pxl_color = 3'b111;
					111	: current_pxl_color = 3'b111;
					112	: current_pxl_color = 3'b111;
					113	: current_pxl_color = 3'b111;
					114	: current_pxl_color = 3'b000;
					115	: current_pxl_color = 3'b000;
					116	: current_pxl_color = 3'b111;
					117	: current_pxl_color = 3'b111;
					118	: current_pxl_color = 3'b111;
					119	: current_pxl_color = 3'b110;
					120	: current_pxl_color = 3'b110;
					121	: current_pxl_color = 3'b111;
					122	: current_pxl_color = 3'b111;
					123	: current_pxl_color = 3'b111;
					124	: current_pxl_color = 3'b000;
					125	: current_pxl_color = 3'b000;
					126	: current_pxl_color = 3'b111;
					127	: current_pxl_color = 3'b111;
					128	: current_pxl_color = 3'b111;
					129	: current_pxl_color = 3'b111;
					130	: current_pxl_color = 3'b000;
					131	: current_pxl_color = 3'b000;
					132	: current_pxl_color = 3'b111;
					133	: current_pxl_color = 3'b111;
					134	: current_pxl_color = 3'b111;
					135	: current_pxl_color = 3'b111;
					136	: current_pxl_color = 3'b111;
					137	: current_pxl_color = 3'b111;
					138	: current_pxl_color = 3'b111;
					139	: current_pxl_color = 3'b111;
					140	: current_pxl_color = 3'b000;
					141	: current_pxl_color = 3'b000;
					142	: current_pxl_color = 3'b111;
					143	: current_pxl_color = 3'b111;
					144	: current_pxl_color = 3'b111;
					145	: current_pxl_color = 3'b111;
					146	: current_pxl_color = 3'b000;
					147	: current_pxl_color = 3'b000;
					148	: current_pxl_color = 3'b111;
					149	: current_pxl_color = 3'b111;
					150	: current_pxl_color = 3'b111;
					151	: current_pxl_color = 3'b111;
					152	: current_pxl_color = 3'b111;
					153	: current_pxl_color = 3'b111;
					154	: current_pxl_color = 3'b111;
					155	: current_pxl_color = 3'b111;
					156	: current_pxl_color = 3'b000;
					157	: current_pxl_color = 3'b000;
					158	: current_pxl_color = 3'b111;
					159	: current_pxl_color = 3'b111;
					160	: current_pxl_color = 3'b111;
					161	: current_pxl_color = 3'b111;
					162	: current_pxl_color = 3'b111;
					163	: current_pxl_color = 3'b000;
					164	: current_pxl_color = 3'b000;
					165	: current_pxl_color = 3'b111;
					166	: current_pxl_color = 3'b111;
					167	: current_pxl_color = 3'b111;
					168	: current_pxl_color = 3'b111;
					169	: current_pxl_color = 3'b111;
					170	: current_pxl_color = 3'b111;
					171	: current_pxl_color = 3'b000;
					172	: current_pxl_color = 3'b000;
					173	: current_pxl_color = 3'b111;
					174	: current_pxl_color = 3'b111;
					175	: current_pxl_color = 3'b111;
					176	: current_pxl_color = 3'b111;
					177	: current_pxl_color = 3'b111;
					178	: current_pxl_color = 3'b111;
					179	: current_pxl_color = 3'b111;
					180	: current_pxl_color = 3'b000;
					181	: current_pxl_color = 3'b111;
					182	: current_pxl_color = 3'b111;
					183	: current_pxl_color = 3'b111;
					184	: current_pxl_color = 3'b111;
					185	: current_pxl_color = 3'b111;
					186	: current_pxl_color = 3'b111;
					187	: current_pxl_color = 3'b000;
					188	: current_pxl_color = 3'b111;
					189	: current_pxl_color = 3'b111;
					190	: current_pxl_color = 3'b111;
					191	: current_pxl_color = 3'b111;
					192	: current_pxl_color = 3'b111;
					193	: current_pxl_color = 3'b111;
					194	: current_pxl_color = 3'b111;
					195	: current_pxl_color = 3'b111;
					196	: current_pxl_color = 3'b000;
					197	: current_pxl_color = 3'b111;
					198	: current_pxl_color = 3'b111;
					199	: current_pxl_color = 3'b111;
					200	: current_pxl_color = 3'b111;
					201	: current_pxl_color = 3'b111;
					202	: current_pxl_color = 3'b111;
					203	: current_pxl_color = 3'b000;
					204	: current_pxl_color = 3'b111;
					205	: current_pxl_color = 3'b111;
					206	: current_pxl_color = 3'b111;
					207	: current_pxl_color = 3'b111;
					208	: current_pxl_color = 3'b111;
					209	: current_pxl_color = 3'b111;
					210	: current_pxl_color = 3'b111;
					211	: current_pxl_color = 3'b111;
					212	: current_pxl_color = 3'b111;
					213	: current_pxl_color = 3'b110;
					214	: current_pxl_color = 3'b110;
					215	: current_pxl_color = 3'b000;
					216	: current_pxl_color = 3'b000;
					217	: current_pxl_color = 3'b110;
					218	: current_pxl_color = 3'b110;
					219	: current_pxl_color = 3'b111;
					220	: current_pxl_color = 3'b111;
					221	: current_pxl_color = 3'b111;
					222	: current_pxl_color = 3'b111;
					223	: current_pxl_color = 3'b111;
					224	: current_pxl_color = 3'b111;
					225	: current_pxl_color = 3'b111;
					226	: current_pxl_color = 3'b111;
					227	: current_pxl_color = 3'b111;
					228	: current_pxl_color = 3'b111;
					229	: current_pxl_color = 3'b111;
					230	: current_pxl_color = 3'b111;
					231	: current_pxl_color = 3'b111;
					232	: current_pxl_color = 3'b111;
					233	: current_pxl_color = 3'b111;
					234	: current_pxl_color = 3'b111;
					235	: current_pxl_color = 3'b111;
					236	: current_pxl_color = 3'b111;
					237	: current_pxl_color = 3'b111;
					238	: current_pxl_color = 3'b111;
					239	: current_pxl_color = 3'b111;
					240	: current_pxl_color = 3'b111;
					241	: current_pxl_color = 3'b111;
					242	: current_pxl_color = 3'b111;
					243	: current_pxl_color = 3'b111;
					244	: current_pxl_color = 3'b111;
					245	: current_pxl_color = 3'b111;
					246	: current_pxl_color = 3'b111;
					247	: current_pxl_color = 3'b111;
					248	: current_pxl_color = 3'b111;
					249	: current_pxl_color = 3'b111;
					250	: current_pxl_color = 3'b111;
					251	: current_pxl_color = 3'b111;
					252	: current_pxl_color = 3'b111;
					253	: current_pxl_color = 3'b111;
					254	: current_pxl_color = 3'b111;
					255	: current_pxl_color = 3'b111;
				endcase
			end
		1 :
			begin
				case (pxl_coor)
					0	: current_pxl_color = 3'b111;
					1	: current_pxl_color = 3'b111;
					2	: current_pxl_color = 3'b111;
					3	: current_pxl_color = 3'b111;
					4	: current_pxl_color = 3'b111;
					5	: current_pxl_color = 3'b111;
					6	: current_pxl_color = 3'b111;
					7	: current_pxl_color = 3'b111;
					8	: current_pxl_color = 3'b111;
					9	: current_pxl_color = 3'b111;
					10	: current_pxl_color = 3'b111;
					11	: current_pxl_color = 3'b111;
					12	: current_pxl_color = 3'b111;
					13	: current_pxl_color = 3'b111;
					14	: current_pxl_color = 3'b111;
					15	: current_pxl_color = 3'b111;
					16	: current_pxl_color = 3'b111;
					17	: current_pxl_color = 3'b111;
					18	: current_pxl_color = 3'b111;
					19	: current_pxl_color = 3'b111;
					20	: current_pxl_color = 3'b111;
					21	: current_pxl_color = 3'b111;
					22	: current_pxl_color = 3'b000;
					23	: current_pxl_color = 3'b000;
					24	: current_pxl_color = 3'b000;
					25	: current_pxl_color = 3'b000;
					26	: current_pxl_color = 3'b111;
					27	: current_pxl_color = 3'b111;
					28	: current_pxl_color = 3'b111;
					29	: current_pxl_color = 3'b111;
					30	: current_pxl_color = 3'b111;
					31	: current_pxl_color = 3'b111;
					32	: current_pxl_color = 3'b111;
					33	: current_pxl_color = 3'b111;
					34	: current_pxl_color = 3'b111;
					35	: current_pxl_color = 3'b111;
					36	: current_pxl_color = 3'b111;
					37	: current_pxl_color = 3'b000;
					38	: current_pxl_color = 3'b000;
					39	: current_pxl_color = 3'b000;
					40	: current_pxl_color = 3'b000;
					41	: current_pxl_color = 3'b000;
					42	: current_pxl_color = 3'b000;
					43	: current_pxl_color = 3'b111;
					44	: current_pxl_color = 3'b111;
					45	: current_pxl_color = 3'b111;
					46	: current_pxl_color = 3'b111;
					47	: current_pxl_color = 3'b111;
					48	: current_pxl_color = 3'b111;
					49	: current_pxl_color = 3'b111;
					50	: current_pxl_color = 3'b111;
					51	: current_pxl_color = 3'b111;
					52	: current_pxl_color = 3'b111;
					53	: current_pxl_color = 3'b000;
					54	: current_pxl_color = 3'b111;
					55	: current_pxl_color = 3'b111;
					56	: current_pxl_color = 3'b111;
					57	: current_pxl_color = 3'b111;
					58	: current_pxl_color = 3'b000;
					59	: current_pxl_color = 3'b111;
					60	: current_pxl_color = 3'b111;
					61	: current_pxl_color = 3'b111;
					62	: current_pxl_color = 3'b111;
					63	: current_pxl_color = 3'b111;
					64	: current_pxl_color = 3'b111;
					65	: current_pxl_color = 3'b111;
					66	: current_pxl_color = 3'b111;
					67	: current_pxl_color = 3'b111;
					68	: current_pxl_color = 3'b111;
					69	: current_pxl_color = 3'b000;
					70	: current_pxl_color = 3'b111;
					71	: current_pxl_color = 3'b000;
					72	: current_pxl_color = 3'b111;
					73	: current_pxl_color = 3'b111;
					74	: current_pxl_color = 3'b000;
					75	: current_pxl_color = 3'b111;
					76	: current_pxl_color = 3'b111;
					77	: current_pxl_color = 3'b111;
					78	: current_pxl_color = 3'b111;
					79	: current_pxl_color = 3'b111;
					80	: current_pxl_color = 3'b111;
					81	: current_pxl_color = 3'b111;
					82	: current_pxl_color = 3'b111;
					83	: current_pxl_color = 3'b111;
					84	: current_pxl_color = 3'b111;
					85	: current_pxl_color = 3'b000;
					86	: current_pxl_color = 3'b111;
					87	: current_pxl_color = 3'b000;
					88	: current_pxl_color = 3'b111;
					89	: current_pxl_color = 3'b111;
					90	: current_pxl_color = 3'b000;
					91	: current_pxl_color = 3'b111;
					92	: current_pxl_color = 3'b111;
					93	: current_pxl_color = 3'b111;
					94	: current_pxl_color = 3'b111;
					95	: current_pxl_color = 3'b111;
					96	: current_pxl_color = 3'b111;
					97	: current_pxl_color = 3'b111;
					98	: current_pxl_color = 3'b111;
					99	: current_pxl_color = 3'b111;
					100	: current_pxl_color = 3'b110;
					101	: current_pxl_color = 3'b110;
					102	: current_pxl_color = 3'b111;
					103	: current_pxl_color = 3'b111;
					104	: current_pxl_color = 3'b111;
					105	: current_pxl_color = 3'b111;
					106	: current_pxl_color = 3'b000;
					107	: current_pxl_color = 3'b111;
					108	: current_pxl_color = 3'b111;
					109	: current_pxl_color = 3'b111;
					110	: current_pxl_color = 3'b111;
					111	: current_pxl_color = 3'b111;
					112	: current_pxl_color = 3'b111;
					113	: current_pxl_color = 3'b111;
					114	: current_pxl_color = 3'b111;
					115	: current_pxl_color = 3'b111;
					116	: current_pxl_color = 3'b111;
					117	: current_pxl_color = 3'b000;
					118	: current_pxl_color = 3'b111;
					119	: current_pxl_color = 3'b000;
					120	: current_pxl_color = 3'b000;
					121	: current_pxl_color = 3'b000;
					122	: current_pxl_color = 3'b000;
					123	: current_pxl_color = 3'b111;
					124	: current_pxl_color = 3'b111;
					125	: current_pxl_color = 3'b111;
					126	: current_pxl_color = 3'b111;
					127	: current_pxl_color = 3'b111;
					128	: current_pxl_color = 3'b111;
					129	: current_pxl_color = 3'b111;
					130	: current_pxl_color = 3'b111;
					131	: current_pxl_color = 3'b111;
					132	: current_pxl_color = 3'b111;
					133	: current_pxl_color = 3'b000;
					134	: current_pxl_color = 3'b111;
					135	: current_pxl_color = 3'b000;
					136	: current_pxl_color = 3'b000;
					137	: current_pxl_color = 3'b000;
					138	: current_pxl_color = 3'b111;
					139	: current_pxl_color = 3'b111;
					140	: current_pxl_color = 3'b111;
					141	: current_pxl_color = 3'b111;
					142	: current_pxl_color = 3'b111;
					143	: current_pxl_color = 3'b111;
					144	: current_pxl_color = 3'b111;
					145	: current_pxl_color = 3'b111;
					146	: current_pxl_color = 3'b111;
					147	: current_pxl_color = 3'b111;
					148	: current_pxl_color = 3'b111;
					149	: current_pxl_color = 3'b000;
					150	: current_pxl_color = 3'b111;
					151	: current_pxl_color = 3'b000;
					152	: current_pxl_color = 3'b000;
					153	: current_pxl_color = 3'b000;
					154	: current_pxl_color = 3'b111;
					155	: current_pxl_color = 3'b111;
					156	: current_pxl_color = 3'b111;
					157	: current_pxl_color = 3'b111;
					158	: current_pxl_color = 3'b111;
					159	: current_pxl_color = 3'b111;
					160	: current_pxl_color = 3'b111;
					161	: current_pxl_color = 3'b111;
					162	: current_pxl_color = 3'b111;
					163	: current_pxl_color = 3'b111;
					164	: current_pxl_color = 3'b111;
					165	: current_pxl_color = 3'b000;
					166	: current_pxl_color = 3'b111;
					167	: current_pxl_color = 3'b000;
					168	: current_pxl_color = 3'b111;
					169	: current_pxl_color = 3'b000;
					170	: current_pxl_color = 3'b111;
					171	: current_pxl_color = 3'b111;
					172	: current_pxl_color = 3'b111;
					173	: current_pxl_color = 3'b111;
					174	: current_pxl_color = 3'b111;
					175	: current_pxl_color = 3'b111;
					176	: current_pxl_color = 3'b111;
					177	: current_pxl_color = 3'b111;
					178	: current_pxl_color = 3'b111;
					179	: current_pxl_color = 3'b111;
					180	: current_pxl_color = 3'b111;
					181	: current_pxl_color = 3'b000;
					182	: current_pxl_color = 3'b111;
					183	: current_pxl_color = 3'b111;
					184	: current_pxl_color = 3'b111;
					185	: current_pxl_color = 3'b000;
					186	: current_pxl_color = 3'b111;
					187	: current_pxl_color = 3'b111;
					188	: current_pxl_color = 3'b111;
					189	: current_pxl_color = 3'b111;
					190	: current_pxl_color = 3'b111;
					191	: current_pxl_color = 3'b111;
					192	: current_pxl_color = 3'b111;
					193	: current_pxl_color = 3'b111;
					194	: current_pxl_color = 3'b111;
					195	: current_pxl_color = 3'b111;
					196	: current_pxl_color = 3'b111;
					197	: current_pxl_color = 3'b000;
					198	: current_pxl_color = 3'b111;
					199	: current_pxl_color = 3'b111;
					200	: current_pxl_color = 3'b000;
					201	: current_pxl_color = 3'b000;
					202	: current_pxl_color = 3'b111;
					203	: current_pxl_color = 3'b111;
					204	: current_pxl_color = 3'b111;
					205	: current_pxl_color = 3'b111;
					206	: current_pxl_color = 3'b111;
					207	: current_pxl_color = 3'b111;
					208	: current_pxl_color = 3'b111;
					209	: current_pxl_color = 3'b111;
					210	: current_pxl_color = 3'b111;
					211	: current_pxl_color = 3'b111;
					212	: current_pxl_color = 3'b110;
					213	: current_pxl_color = 3'b110;
					214	: current_pxl_color = 3'b000;
					215	: current_pxl_color = 3'b000;
					216	: current_pxl_color = 3'b000;
					217	: current_pxl_color = 3'b111;
					218	: current_pxl_color = 3'b111;
					219	: current_pxl_color = 3'b111;
					220	: current_pxl_color = 3'b111;
					221	: current_pxl_color = 3'b111;
					222	: current_pxl_color = 3'b111;
					223	: current_pxl_color = 3'b111;
					224	: current_pxl_color = 3'b111;
					225	: current_pxl_color = 3'b111;
					226	: current_pxl_color = 3'b111;
					227	: current_pxl_color = 3'b111;
					228	: current_pxl_color = 3'b111;
					229	: current_pxl_color = 3'b111;
					230	: current_pxl_color = 3'b111;
					231	: current_pxl_color = 3'b111;
					232	: current_pxl_color = 3'b111;
					233	: current_pxl_color = 3'b111;
					234	: current_pxl_color = 3'b111;
					235	: current_pxl_color = 3'b111;
					236	: current_pxl_color = 3'b111;
					237	: current_pxl_color = 3'b111;
					238	: current_pxl_color = 3'b111;
					239	: current_pxl_color = 3'b111;
					240	: current_pxl_color = 3'b111;
					241	: current_pxl_color = 3'b111;
					242	: current_pxl_color = 3'b111;
					243	: current_pxl_color = 3'b111;
					244	: current_pxl_color = 3'b111;
					245	: current_pxl_color = 3'b111;
					246	: current_pxl_color = 3'b111;
					247	: current_pxl_color = 3'b111;
					248	: current_pxl_color = 3'b111;
					249	: current_pxl_color = 3'b111;
					250	: current_pxl_color = 3'b111;
					251	: current_pxl_color = 3'b111;
					252	: current_pxl_color = 3'b111;
					253	: current_pxl_color = 3'b111;
					254	: current_pxl_color = 3'b111;
					255	: current_pxl_color = 3'b111;
				endcase
			end
		3 :
			begin
				case (pxl_coor)
					0	: current_pxl_color = 3'b111;
					1	: current_pxl_color = 3'b111;
					2	: current_pxl_color = 3'b111;
					3	: current_pxl_color = 3'b111;
					4	: current_pxl_color = 3'b111;
					5	: current_pxl_color = 3'b111;
					6	: current_pxl_color = 3'b111;
					7	: current_pxl_color = 3'b111;
					8	: current_pxl_color = 3'b111;
					9	: current_pxl_color = 3'b111;
					10	: current_pxl_color = 3'b111;
					11	: current_pxl_color = 3'b111;
					12	: current_pxl_color = 3'b111;
					13	: current_pxl_color = 3'b111;
					14	: current_pxl_color = 3'b111;
					15	: current_pxl_color = 3'b111;
					16	: current_pxl_color = 3'b111;
					17	: current_pxl_color = 3'b111;
					18	: current_pxl_color = 3'b111;
					19	: current_pxl_color = 3'b111;
					20	: current_pxl_color = 3'b111;
					21	: current_pxl_color = 3'b111;
					22	: current_pxl_color = 3'b000;
					23	: current_pxl_color = 3'b000;
					24	: current_pxl_color = 3'b000;
					25	: current_pxl_color = 3'b000;
					26	: current_pxl_color = 3'b111;
					27	: current_pxl_color = 3'b111;
					28	: current_pxl_color = 3'b111;
					29	: current_pxl_color = 3'b111;
					30	: current_pxl_color = 3'b111;
					31	: current_pxl_color = 3'b111;
					32	: current_pxl_color = 3'b111;
					33	: current_pxl_color = 3'b111;
					34	: current_pxl_color = 3'b111;
					35	: current_pxl_color = 3'b111;
					36	: current_pxl_color = 3'b111;
					37	: current_pxl_color = 3'b000;
					38	: current_pxl_color = 3'b000;
					39	: current_pxl_color = 3'b111;
					40	: current_pxl_color = 3'b111;
					41	: current_pxl_color = 3'b000;
					42	: current_pxl_color = 3'b000;
					43	: current_pxl_color = 3'b111;
					44	: current_pxl_color = 3'b111;
					45	: current_pxl_color = 3'b111;
					46	: current_pxl_color = 3'b111;
					47	: current_pxl_color = 3'b111;
					48	: current_pxl_color = 3'b111;
					49	: current_pxl_color = 3'b111;
					50	: current_pxl_color = 3'b111;
					51	: current_pxl_color = 3'b111;
					52	: current_pxl_color = 3'b111;
					53	: current_pxl_color = 3'b000;
					54	: current_pxl_color = 3'b111;
					55	: current_pxl_color = 3'b111;
					56	: current_pxl_color = 3'b111;
					57	: current_pxl_color = 3'b111;
					58	: current_pxl_color = 3'b000;
					59	: current_pxl_color = 3'b111;
					60	: current_pxl_color = 3'b111;
					61	: current_pxl_color = 3'b111;
					62	: current_pxl_color = 3'b111;
					63	: current_pxl_color = 3'b111;
					64	: current_pxl_color = 3'b111;
					65	: current_pxl_color = 3'b111;
					66	: current_pxl_color = 3'b111;
					67	: current_pxl_color = 3'b111;
					68	: current_pxl_color = 3'b111;
					69	: current_pxl_color = 3'b000;
					70	: current_pxl_color = 3'b111;
					71	: current_pxl_color = 3'b111;
					72	: current_pxl_color = 3'b000;
					73	: current_pxl_color = 3'b111;
					74	: current_pxl_color = 3'b000;
					75	: current_pxl_color = 3'b111;
					76	: current_pxl_color = 3'b111;
					77	: current_pxl_color = 3'b111;
					78	: current_pxl_color = 3'b111;
					79	: current_pxl_color = 3'b111;
					80	: current_pxl_color = 3'b111;
					81	: current_pxl_color = 3'b111;
					82	: current_pxl_color = 3'b111;
					83	: current_pxl_color = 3'b111;
					84	: current_pxl_color = 3'b111;
					85	: current_pxl_color = 3'b000;
					86	: current_pxl_color = 3'b111;
					87	: current_pxl_color = 3'b111;
					88	: current_pxl_color = 3'b000;
					89	: current_pxl_color = 3'b111;
					90	: current_pxl_color = 3'b000;
					91	: current_pxl_color = 3'b111;
					92	: current_pxl_color = 3'b111;
					93	: current_pxl_color = 3'b111;
					94	: current_pxl_color = 3'b111;
					95	: current_pxl_color = 3'b111;
					96	: current_pxl_color = 3'b111;
					97	: current_pxl_color = 3'b111;
					98	: current_pxl_color = 3'b111;
					99	: current_pxl_color = 3'b111;
					100	: current_pxl_color = 3'b111;
					101	: current_pxl_color = 3'b000;
					102	: current_pxl_color = 3'b111;
					103	: current_pxl_color = 3'b111;
					104	: current_pxl_color = 3'b111;
					105	: current_pxl_color = 3'b111;
					106	: current_pxl_color = 3'b110;
					107	: current_pxl_color = 3'b110;
					108	: current_pxl_color = 3'b111;
					109	: current_pxl_color = 3'b111;
					110	: current_pxl_color = 3'b111;
					111	: current_pxl_color = 3'b111;
					112	: current_pxl_color = 3'b111;
					113	: current_pxl_color = 3'b111;
					114	: current_pxl_color = 3'b111;
					115	: current_pxl_color = 3'b111;
					116	: current_pxl_color = 3'b111;
					117	: current_pxl_color = 3'b000;
					118	: current_pxl_color = 3'b000;
					119	: current_pxl_color = 3'b000;
					120	: current_pxl_color = 3'b000;
					121	: current_pxl_color = 3'b111;
					122	: current_pxl_color = 3'b000;
					123	: current_pxl_color = 3'b111;
					124	: current_pxl_color = 3'b111;
					125	: current_pxl_color = 3'b111;
					126	: current_pxl_color = 3'b111;
					127	: current_pxl_color = 3'b111;
					128	: current_pxl_color = 3'b111;
					129	: current_pxl_color = 3'b111;
					130	: current_pxl_color = 3'b111;
					131	: current_pxl_color = 3'b111;
					132	: current_pxl_color = 3'b111;
					133	: current_pxl_color = 3'b111;
					134	: current_pxl_color = 3'b000;
					135	: current_pxl_color = 3'b000;
					136	: current_pxl_color = 3'b000;
					137	: current_pxl_color = 3'b111;
					138	: current_pxl_color = 3'b000;
					139	: current_pxl_color = 3'b111;
					140	: current_pxl_color = 3'b111;
					141	: current_pxl_color = 3'b111;
					142	: current_pxl_color = 3'b111;
					143	: current_pxl_color = 3'b111;
					144	: current_pxl_color = 3'b111;
					145	: current_pxl_color = 3'b111;
					146	: current_pxl_color = 3'b111;
					147	: current_pxl_color = 3'b111;
					148	: current_pxl_color = 3'b111;
					149	: current_pxl_color = 3'b111;
					150	: current_pxl_color = 3'b000;
					151	: current_pxl_color = 3'b000;
					152	: current_pxl_color = 3'b000;
					153	: current_pxl_color = 3'b111;
					154	: current_pxl_color = 3'b000;
					155	: current_pxl_color = 3'b111;
					156	: current_pxl_color = 3'b111;
					157	: current_pxl_color = 3'b111;
					158	: current_pxl_color = 3'b111;
					159	: current_pxl_color = 3'b111;
					160	: current_pxl_color = 3'b111;
					161	: current_pxl_color = 3'b111;
					162	: current_pxl_color = 3'b111;
					163	: current_pxl_color = 3'b111;
					164	: current_pxl_color = 3'b111;
					165	: current_pxl_color = 3'b111;
					166	: current_pxl_color = 3'b000;
					167	: current_pxl_color = 3'b111;
					168	: current_pxl_color = 3'b000;
					169	: current_pxl_color = 3'b111;
					170	: current_pxl_color = 3'b000;
					171	: current_pxl_color = 3'b111;
					172	: current_pxl_color = 3'b111;
					173	: current_pxl_color = 3'b111;
					174	: current_pxl_color = 3'b111;
					175	: current_pxl_color = 3'b111;
					176	: current_pxl_color = 3'b111;
					177	: current_pxl_color = 3'b111;
					178	: current_pxl_color = 3'b111;
					179	: current_pxl_color = 3'b111;
					180	: current_pxl_color = 3'b111;
					181	: current_pxl_color = 3'b111;
					182	: current_pxl_color = 3'b000;
					183	: current_pxl_color = 3'b111;
					184	: current_pxl_color = 3'b111;
					185	: current_pxl_color = 3'b111;
					186	: current_pxl_color = 3'b000;
					187	: current_pxl_color = 3'b111;
					188	: current_pxl_color = 3'b111;
					189	: current_pxl_color = 3'b111;
					190	: current_pxl_color = 3'b111;
					191	: current_pxl_color = 3'b111;
					192	: current_pxl_color = 3'b111;
					193	: current_pxl_color = 3'b111;
					194	: current_pxl_color = 3'b111;
					195	: current_pxl_color = 3'b111;
					196	: current_pxl_color = 3'b111;
					197	: current_pxl_color = 3'b111;
					198	: current_pxl_color = 3'b000;
					199	: current_pxl_color = 3'b000;
					200	: current_pxl_color = 3'b111;
					201	: current_pxl_color = 3'b111;
					202	: current_pxl_color = 3'b000;
					203	: current_pxl_color = 3'b111;
					204	: current_pxl_color = 3'b111;
					205	: current_pxl_color = 3'b111;
					206	: current_pxl_color = 3'b111;
					207	: current_pxl_color = 3'b111;
					208	: current_pxl_color = 3'b111;
					209	: current_pxl_color = 3'b111;
					210	: current_pxl_color = 3'b111;
					211	: current_pxl_color = 3'b111;
					212	: current_pxl_color = 3'b111;
					213	: current_pxl_color = 3'b111;
					214	: current_pxl_color = 3'b111;
					215	: current_pxl_color = 3'b000;
					216	: current_pxl_color = 3'b000;
					217	: current_pxl_color = 3'b000;
					218	: current_pxl_color = 3'b110;
					219	: current_pxl_color = 3'b110;
					220	: current_pxl_color = 3'b111;
					221	: current_pxl_color = 3'b111;
					222	: current_pxl_color = 3'b111;
					223	: current_pxl_color = 3'b111;
					224	: current_pxl_color = 3'b111;
					225	: current_pxl_color = 3'b111;
					226	: current_pxl_color = 3'b111;
					227	: current_pxl_color = 3'b111;
					228	: current_pxl_color = 3'b111;
					229	: current_pxl_color = 3'b111;
					230	: current_pxl_color = 3'b111;
					231	: current_pxl_color = 3'b111;
					232	: current_pxl_color = 3'b111;
					233	: current_pxl_color = 3'b111;
					234	: current_pxl_color = 3'b111;
					235	: current_pxl_color = 3'b111;
					236	: current_pxl_color = 3'b111;
					237	: current_pxl_color = 3'b111;
					238	: current_pxl_color = 3'b111;
					239	: current_pxl_color = 3'b111;
					240	: current_pxl_color = 3'b111;
					241	: current_pxl_color = 3'b111;
					242	: current_pxl_color = 3'b111;
					243	: current_pxl_color = 3'b111;
					244	: current_pxl_color = 3'b111;
					245	: current_pxl_color = 3'b111;
					246	: current_pxl_color = 3'b111;
					247	: current_pxl_color = 3'b111;
					248	: current_pxl_color = 3'b111;
					249	: current_pxl_color = 3'b111;
					250	: current_pxl_color = 3'b111;
					251	: current_pxl_color = 3'b111;
					252	: current_pxl_color = 3'b111;
					253	: current_pxl_color = 3'b111;
					254	: current_pxl_color = 3'b111;
					255	: current_pxl_color = 3'b111;
				endcase
			end
		2 :
			begin
				case (pxl_coor)
					0	: current_pxl_color = 3'b111;
					1	: current_pxl_color = 3'b111;
					2	: current_pxl_color = 3'b111;
					3	: current_pxl_color = 3'b111;
					4	: current_pxl_color = 3'b111;
					5	: current_pxl_color = 3'b111;
					6	: current_pxl_color = 3'b111;
					7	: current_pxl_color = 3'b111;
					8	: current_pxl_color = 3'b111;
					9	: current_pxl_color = 3'b111;
					10	: current_pxl_color = 3'b111;
					11	: current_pxl_color = 3'b111;
					12	: current_pxl_color = 3'b111;
					13	: current_pxl_color = 3'b111;
					14	: current_pxl_color = 3'b111;
					15	: current_pxl_color = 3'b111;
					16	: current_pxl_color = 3'b111;
					17	: current_pxl_color = 3'b111;
					18	: current_pxl_color = 3'b111;
					19	: current_pxl_color = 3'b111;
					20	: current_pxl_color = 3'b111;
					21	: current_pxl_color = 3'b111;
					22	: current_pxl_color = 3'b000;
					23	: current_pxl_color = 3'b000;
					24	: current_pxl_color = 3'b000;
					25	: current_pxl_color = 3'b000;
					26	: current_pxl_color = 3'b111;
					27	: current_pxl_color = 3'b111;
					28	: current_pxl_color = 3'b111;
					29	: current_pxl_color = 3'b111;
					30	: current_pxl_color = 3'b111;
					31	: current_pxl_color = 3'b111;
					32	: current_pxl_color = 3'b111;
					33	: current_pxl_color = 3'b111;
					34	: current_pxl_color = 3'b111;
					35	: current_pxl_color = 3'b111;
					36	: current_pxl_color = 3'b111;
					37	: current_pxl_color = 3'b000;
					38	: current_pxl_color = 3'b000;
					39	: current_pxl_color = 3'b000;
					40	: current_pxl_color = 3'b000;
					41	: current_pxl_color = 3'b000;
					42	: current_pxl_color = 3'b000;
					43	: current_pxl_color = 3'b111;
					44	: current_pxl_color = 3'b111;
					45	: current_pxl_color = 3'b111;
					46	: current_pxl_color = 3'b111;
					47	: current_pxl_color = 3'b111;
					48	: current_pxl_color = 3'b111;
					49	: current_pxl_color = 3'b111;
					50	: current_pxl_color = 3'b111;
					51	: current_pxl_color = 3'b111;
					52	: current_pxl_color = 3'b000;
					53	: current_pxl_color = 3'b000;
					54	: current_pxl_color = 3'b000;
					55	: current_pxl_color = 3'b000;
					56	: current_pxl_color = 3'b000;
					57	: current_pxl_color = 3'b000;
					58	: current_pxl_color = 3'b000;
					59	: current_pxl_color = 3'b000;
					60	: current_pxl_color = 3'b111;
					61	: current_pxl_color = 3'b111;
					62	: current_pxl_color = 3'b111;
					63	: current_pxl_color = 3'b111;
					64	: current_pxl_color = 3'b111;
					65	: current_pxl_color = 3'b111;
					66	: current_pxl_color = 3'b111;
					67	: current_pxl_color = 3'b111;
					68	: current_pxl_color = 3'b000;
					69	: current_pxl_color = 3'b000;
					70	: current_pxl_color = 3'b000;
					71	: current_pxl_color = 3'b000;
					72	: current_pxl_color = 3'b000;
					73	: current_pxl_color = 3'b000;
					74	: current_pxl_color = 3'b000;
					75	: current_pxl_color = 3'b000;
					76	: current_pxl_color = 3'b111;
					77	: current_pxl_color = 3'b111;
					78	: current_pxl_color = 3'b111;
					79	: current_pxl_color = 3'b111;
					80	: current_pxl_color = 3'b111;
					81	: current_pxl_color = 3'b111;
					82	: current_pxl_color = 3'b111;
					83	: current_pxl_color = 3'b111;
					84	: current_pxl_color = 3'b000;
					85	: current_pxl_color = 3'b000;
					86	: current_pxl_color = 3'b000;
					87	: current_pxl_color = 3'b000;
					88	: current_pxl_color = 3'b000;
					89	: current_pxl_color = 3'b000;
					90	: current_pxl_color = 3'b000;
					91	: current_pxl_color = 3'b000;
					92	: current_pxl_color = 3'b111;
					93	: current_pxl_color = 3'b111;
					94	: current_pxl_color = 3'b111;
					95	: current_pxl_color = 3'b111;
					96	: current_pxl_color = 3'b111;
					97	: current_pxl_color = 3'b111;
					98	: current_pxl_color = 3'b111;
					99	: current_pxl_color = 3'b000;
					100	: current_pxl_color = 3'b000;
					101	: current_pxl_color = 3'b000;
					102	: current_pxl_color = 3'b000;
					103	: current_pxl_color = 3'b000;
					104	: current_pxl_color = 3'b000;
					105	: current_pxl_color = 3'b000;
					106	: current_pxl_color = 3'b000;
					107	: current_pxl_color = 3'b000;
					108	: current_pxl_color = 3'b000;
					109	: current_pxl_color = 3'b111;
					110	: current_pxl_color = 3'b111;
					111	: current_pxl_color = 3'b111;
					112	: current_pxl_color = 3'b111;
					113	: current_pxl_color = 3'b111;
					114	: current_pxl_color = 3'b000;
					115	: current_pxl_color = 3'b000;
					116	: current_pxl_color = 3'b000;
					117	: current_pxl_color = 3'b000;
					118	: current_pxl_color = 3'b000;
					119	: current_pxl_color = 3'b000;
					120	: current_pxl_color = 3'b000;
					121	: current_pxl_color = 3'b000;
					122	: current_pxl_color = 3'b000;
					123	: current_pxl_color = 3'b000;
					124	: current_pxl_color = 3'b000;
					125	: current_pxl_color = 3'b000;
					126	: current_pxl_color = 3'b111;
					127	: current_pxl_color = 3'b111;
					128	: current_pxl_color = 3'b111;
					129	: current_pxl_color = 3'b111;
					130	: current_pxl_color = 3'b000;
					131	: current_pxl_color = 3'b000;
					132	: current_pxl_color = 3'b000;
					133	: current_pxl_color = 3'b000;
					134	: current_pxl_color = 3'b000;
					135	: current_pxl_color = 3'b000;
					136	: current_pxl_color = 3'b000;
					137	: current_pxl_color = 3'b000;
					138	: current_pxl_color = 3'b000;
					139	: current_pxl_color = 3'b000;
					140	: current_pxl_color = 3'b000;
					141	: current_pxl_color = 3'b000;
					142	: current_pxl_color = 3'b111;
					143	: current_pxl_color = 3'b111;
					144	: current_pxl_color = 3'b111;
					145	: current_pxl_color = 3'b111;
					146	: current_pxl_color = 3'b000;
					147	: current_pxl_color = 3'b111;
					148	: current_pxl_color = 3'b000;
					149	: current_pxl_color = 3'b000;
					150	: current_pxl_color = 3'b000;
					151	: current_pxl_color = 3'b000;
					152	: current_pxl_color = 3'b000;
					153	: current_pxl_color = 3'b000;
					154	: current_pxl_color = 3'b000;
					155	: current_pxl_color = 3'b000;
					156	: current_pxl_color = 3'b111;
					157	: current_pxl_color = 3'b000;
					158	: current_pxl_color = 3'b111;
					159	: current_pxl_color = 3'b111;
					160	: current_pxl_color = 3'b111;
					161	: current_pxl_color = 3'b111;
					162	: current_pxl_color = 3'b111;
					163	: current_pxl_color = 3'b111;
					164	: current_pxl_color = 3'b000;
					165	: current_pxl_color = 3'b000;
					166	: current_pxl_color = 3'b000;
					167	: current_pxl_color = 3'b000;
					168	: current_pxl_color = 3'b000;
					169	: current_pxl_color = 3'b000;
					170	: current_pxl_color = 3'b000;
					171	: current_pxl_color = 3'b000;
					172	: current_pxl_color = 3'b111;
					173	: current_pxl_color = 3'b111;
					174	: current_pxl_color = 3'b111;
					175	: current_pxl_color = 3'b111;
					176	: current_pxl_color = 3'b111;
					177	: current_pxl_color = 3'b111;
					178	: current_pxl_color = 3'b111;
					179	: current_pxl_color = 3'b111;
					180	: current_pxl_color = 3'b000;
					181	: current_pxl_color = 3'b000;
					182	: current_pxl_color = 3'b000;
					183	: current_pxl_color = 3'b000;
					184	: current_pxl_color = 3'b000;
					185	: current_pxl_color = 3'b000;
					186	: current_pxl_color = 3'b000;
					187	: current_pxl_color = 3'b000;
					188	: current_pxl_color = 3'b111;
					189	: current_pxl_color = 3'b111;
					190	: current_pxl_color = 3'b111;
					191	: current_pxl_color = 3'b111;
					192	: current_pxl_color = 3'b111;
					193	: current_pxl_color = 3'b111;
					194	: current_pxl_color = 3'b111;
					195	: current_pxl_color = 3'b111;
					196	: current_pxl_color = 3'b000;
					197	: current_pxl_color = 3'b000;
					198	: current_pxl_color = 3'b000;
					199	: current_pxl_color = 3'b000;
					200	: current_pxl_color = 3'b000;
					201	: current_pxl_color = 3'b000;
					202	: current_pxl_color = 3'b000;
					203	: current_pxl_color = 3'b000;
					204	: current_pxl_color = 3'b111;
					205	: current_pxl_color = 3'b111;
					206	: current_pxl_color = 3'b111;
					207	: current_pxl_color = 3'b111;
					208	: current_pxl_color = 3'b111;
					209	: current_pxl_color = 3'b111;
					210	: current_pxl_color = 3'b111;
					211	: current_pxl_color = 3'b111;
					212	: current_pxl_color = 3'b111;
					213	: current_pxl_color = 3'b110;
					214	: current_pxl_color = 3'b110;
					215	: current_pxl_color = 3'b000;
					216	: current_pxl_color = 3'b000;
					217	: current_pxl_color = 3'b110;
					218	: current_pxl_color = 3'b110;
					219	: current_pxl_color = 3'b111;
					220	: current_pxl_color = 3'b111;
					221	: current_pxl_color = 3'b111;
					222	: current_pxl_color = 3'b111;
					223	: current_pxl_color = 3'b111;
					224	: current_pxl_color = 3'b111;
					225	: current_pxl_color = 3'b111;
					226	: current_pxl_color = 3'b111;
					227	: current_pxl_color = 3'b111;
					228	: current_pxl_color = 3'b111;
					229	: current_pxl_color = 3'b111;
					230	: current_pxl_color = 3'b111;
					231	: current_pxl_color = 3'b111;
					232	: current_pxl_color = 3'b111;
					233	: current_pxl_color = 3'b111;
					234	: current_pxl_color = 3'b111;
					235	: current_pxl_color = 3'b111;
					236	: current_pxl_color = 3'b111;
					237	: current_pxl_color = 3'b111;
					238	: current_pxl_color = 3'b111;
					239	: current_pxl_color = 3'b111;
					240	: current_pxl_color = 3'b111;
					241	: current_pxl_color = 3'b111;
					242	: current_pxl_color = 3'b111;
					243	: current_pxl_color = 3'b111;
					244	: current_pxl_color = 3'b111;
					245	: current_pxl_color = 3'b111;
					246	: current_pxl_color = 3'b111;
					247	: current_pxl_color = 3'b111;
					248	: current_pxl_color = 3'b111;
					249	: current_pxl_color = 3'b111;
					250	: current_pxl_color = 3'b111;
					251	: current_pxl_color = 3'b111;
					252	: current_pxl_color = 3'b111;
					253	: current_pxl_color = 3'b111;
					254	: current_pxl_color = 3'b111;
					255	: current_pxl_color = 3'b111;
            endcase
        end
	
	endcase
end

assign color = current_pxl_color;

endmodule

